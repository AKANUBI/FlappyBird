//-------------------------------------------------------------------------
//      stair.sv                                                         --
//      Created by Yuhao Ge & Haina Lou                                  --
//      Fall 2021                                                        --
//                                                                       --
//      This module is used to generate stairs                           --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------

// NIO-2 give messages to control the status of the stairs
// The new positon is ramdomlly generated by NOI-2

module pipe ( input Clk, Reset,
					input frame_clk,  
					input [19:0]  random_num,
					input [9:0]   DrawX, DrawY,       
					input [1:0] game_state,
					output logic  is_pipe, is_pipe_edge, is_grd_y, is_grd_g_d, is_grd_g_l,
					output logic [18:0] p_addr, p_e_addr,
					output logic [6:0] score1
					);	                                                                                                                                                                                
					
	 parameter [9:0] width = 10'd50;
	 parameter [9:0] height = 10'd480;
	 parameter [9:0] pipe_X_corner1 = 10'd480;  // left up corner of the pipe
	 parameter [9:0] pipe_X_corner2 = 10'd665;  // left up corner of the pipe
    parameter [9:0] pipe_Y_corner = 10'd0;  // left up corner of the pipe

    
    logic [9:0] pipe_X_Pos1, pipe_X_Pos2, pipe_Y_Pos;
    logic [9:0] pipe_X_Pos_in1, pipe_X_Pos_in2;
	 logic [9:0] bg_pos, bg_pos_in;
	 logic [9:0] random_number1, random_number2, random1_in, random2_in;
	 logic [9:0] random1, random2;
	 logic [6:0] score1_in;
//	 int r,r_in;
//	 logic clk_out;
    //////// Do not modify the always_ff blocks. ////////
    // Detect rising edge of frame_clk
    logic frame_clk_delayed, frame_clk_rising_edge;
    always_ff @ (posedge Clk) begin
        frame_clk_delayed <= frame_clk;
        frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
    end
    // Update registers
	 // Default period (in time units) for the clock
		// Default period (in time units) for the clock
//		parameter PERIOD = 2000000000; // Change this value to set the clock period
//
//		// Internal state variable to keep track of the clock
//		logic state = 0;
//
//		// Clock generation process
//		always @(posedge Clk) begin
//			 #(PERIOD); // Delay for of the clock period
//			 state <= ~state; // Toggle the state
//			 clk_out <= state;
//		end

		// Assign the generated clock to the output port
	 initial begin
      pipe_X_Pos1 <= pipe_X_corner1;
		pipe_X_Pos2 <= pipe_X_corner2;
		pipe_Y_Pos <= pipe_Y_corner;
		bg_pos <= bg_pos_in;
		random1 <= random_num;
		random2 <= random_num-50;
		score1 <= 0;
    end
	 
    always_ff @ (posedge Clk)
    begin
        if (Reset)
        begin
            pipe_X_Pos1 <= pipe_X_corner1;
				pipe_X_Pos2 <= pipe_X_corner2;
				pipe_Y_Pos <= pipe_Y_corner;
				bg_pos <= pipe_X_corner1;
				random1 <= random_num;
				random2 <= random_num-50;
				score1 <= 0;
//				r <= 8'b11111111;
				//pipe_Y_Step <= 10'd1;
        end
        else
        begin
            pipe_X_Pos1 <= pipe_X_Pos_in1;
				pipe_X_Pos2 <= pipe_X_Pos_in2;
				
				score1 <= score1_in;
				
				bg_pos <= bg_pos_in;
				
				random1 <= random1_in;
				random2 <= random2_in;
        end
		  
    end
    //////// Do not modify the always_ff blocks. ////////
	 
//	LFSR rand_num_instance1(.Clk(frame_clk), .r(r), .random_number(random_number1));
//	LFSR rand_num_instance2(.Clk(frame_clk), .random_number(random_number2));  

			
    always_comb
		begin
			pipe_X_Pos_in1 = pipe_X_Pos1;
			pipe_X_Pos_in2 = pipe_X_Pos2;
			bg_pos_in = bg_pos;
			random1_in = random1;
			random2_in = random2;
			score1_in =score1;
	 
			   if (frame_clk_rising_edge) begin

						case (game_state)
							2'd2: begin
								bg_pos_in = bg_pos;
							end
							default: begin
								if (bg_pos <= 10'd160) begin
									bg_pos_in = pipe_X_corner1;
								end else begin
									bg_pos_in = bg_pos - 10'd1;
								end
							end
						endcase
					
					
					case (game_state)
						 2'd1: begin
						 if (pipe_X_Pos1<= 10'd100) begin
							random1_in = random_num;
							pipe_X_Pos_in1 = pipe_X_corner1;
						 end else begin
							  pipe_X_Pos_in1 = pipe_X_Pos1 - 10'd1;
							  if(pipe_X_Pos1 == 290) begin
									score1_in = score1+1;
								end
						 end
						 
						 if (pipe_X_Pos2<= 10'd100) begin
							random2_in = random_num;
							pipe_X_Pos_in2 = pipe_X_corner1;
						 end else begin
							  pipe_X_Pos_in2 = pipe_X_Pos2 - 10'd1;
							  if(pipe_X_Pos2 == 290) begin
									score1_in = score1+1;
								end
						 end
							
						 end

						 2'd2: begin
							  pipe_X_Pos_in1 = pipe_X_Pos1;
							  pipe_X_Pos_in2 = pipe_X_Pos2;
						 end

						 2'd0: begin
							  pipe_X_Pos_in1 = pipe_X_corner1;
							  pipe_X_Pos_in2 = pipe_X_corner2;
							  score1_in = 0;
						 end

						 default: begin
							  pipe_X_Pos_in1 = pipe_X_Pos1;
							  pipe_X_Pos_in2 = pipe_X_Pos2;
						 end
					endcase

						
					
					end
				
				
				
		  end


    // Compute whether the pixel corresponds to pipe or background
    /* Since the multiplicants are required to be signed, we have to first cast them
       from logic to int (signed by default) before they are multiplied. */
    int DistX1, DistX2, DistY, DistX, ran1, ran2;
    assign DistX1 = DrawX - pipe_X_Pos1;
	 assign DistX2 = DrawX - pipe_X_Pos2;
    assign DistY = DrawY - pipe_Y_Pos;
	 assign DistX = DrawX - bg_pos;
	 assign ran1 = random1;
	 assign ran2 = random2;
	 
	 parameter [9:0] width_p_e = 10'd60;

	
    always_comb begin

        if ( (DistX1 < width + 5 && DistX1 >= 5) &&  ((DistY < ran1 - 70 && DistY >= 0)||(DistY >= ran1 + 80 && DistY <= 10'd439))) begin
            is_pipe = 1'b1;
				p_addr = DistX1 - 5;
			end
		else if ( (DistX2 < width +5 && DistX2 >= 5) &&  ((DistY < ran2 - 70 && DistY >= 0)||(DistY >= ran2 + 80 && DistY <= 10'd439))) begin
            is_pipe = 1'b1;
				p_addr = DistX2 - 5;
		  end
        else begin
            is_pipe = 1'b0;
				p_addr = 0;
			end
				
		  if ( (DistX1 < width +10 && DistX1 >= 0) &&  ((DistY <= ran1 - 40 && DistY >= ran1 - 70)||(DistY >= ran1 + 50 && DistY < ran1 + 80))) begin
				is_pipe_edge = 1'b1;
				if (DistY == ran1 - 40 || DistY == ran1 - 70 || DistY == ran1 + 50 || DistY == ran1 + 80) begin
					p_e_addr = DistX1;
				end
				else begin
					p_e_addr = DistX1 + 60;
				end

			end
				
		else if ( (DistX2 < width +10 && DistX2 >= 0) &&  ((DistY <= ran2 - 40 && DistY >= ran2 - 70)||(DistY >= ran2 + 50 && DistY < ran2 + 80))) begin
				is_pipe_edge = 1'b1;
				if (DistY == ran2 - 40 || DistY == ran2 - 70 || DistY == ran2 + 50 || DistY == ran2 + 80) begin
					p_e_addr = DistX2;
				end
				else begin
					p_e_addr = DistX2 + 60;
				end

		end
				
		  else begin
				is_pipe_edge = 1'b0; // pipe edge: 60*10
				p_e_addr = 19'b0;
			end
			
			if (DistY <= 10'd479 && DistY > 10'd444) begin
				is_grd_y = 1'b1;
			end
			else begin
				is_grd_y = 1'b0;
			end
		  
		  if (DistY <= 10'd444 && DistY > 10'd439) begin
				if (DistX < 0 && -DistX % 10 < 5) begin
					is_grd_g_d = 1'b1;
				   is_grd_g_l = 1'b0;
			   end
				
				else if (DistX >= 0 && DistX % 10 >= 5) begin
					is_grd_g_d = 1'b1;
				   is_grd_g_l = 1'b0;
			   end
				
				else begin
					is_grd_g_d = 1'b0;
				   is_grd_g_l = 1'b1;
			   end
			end
			
			else begin
				is_grd_g_d = 1'b0;
				is_grd_g_l = 1'b0;
			end	
        /* The pipe's (pixelated) circle is generated using the standard circle formula.  Note that while 
           the single line is quite powerful descriptively, it causes the synthesis tool to use up three
           of the 12 available multipliers on the chip! */
    end
	 
endmodule